Standard cell Simulation

.include "/home/matt/work/asic-workshop/shuttle2-mpw-two-c/pdk/skywater-pdk/libraries/sky130_fd_pr/latest/models/corners/tt.spice"
.include "top.spice"

Xpoc but_0 but_1 but_2 but_3 but_4 but_5 but_6 but_7 but_8 but_9 clk lock open reset VPWR VGND top
* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

Vbut_0 but_0 VGND 1.8
Vbut_1 but_1 VGND 0
Vbut_2 but_2 VGND 1.8
Vbut_3 but_3 VGND 0
Vbut_4 but_4 VGND 1.8
Vbut_5 but_5 VGND 0
Vbut_6 but_6 VGND 1.8
Vbut_7 but_7 VGND 0
Vbut_8 but_8 VGND 0
Vbut_9 but_9 VGND 0
Vopen open VGND 1.8

*Rlock lock VPWR 10k
* create a clock, 4ns period
* initial v, pulse v, delay, rise, fall, pulse w, period
Vclk clk VGND pulse(0 1.8 1n 10p 10p 2n 4n)

* create reset
* start high, for 4ns, rest of the time off
Vreset reset VGND pulse(0 1.8 0n 10p 10p 2n 20n)

* press the open button
* start low, wait for 4ns, hold high
* Vopen open VGND pulse(0 1.8 4n 10p 10p 20n 20n)

* setup the transient analysis
.tran 10p 20n 0

.control
run
set color0 = white
set color1 = black
plot clk, reset, open, lock
.endc

.end

